`timescale 1ns / 1ps

module pc(input [31:0] i, output reg [31:0] o) ; always @(i) begin o=i; end endmodule
