`timescale 1ns / 1ps


module imem(input clock, input [31:0] addr, output reg [31:0] insto, output reg [31:0] ip, output reg [31:0] idp);
reg [31:0] data [255:0];
initial begin 
//data[0] = 32'b00000000000000000000000000000000;
//data[1] = 32'b00000000000000000000000000000000;
//data[2] = 32'b00110000000000100000110000000000;
//data[3] = 32'b11101000000000100000000000000000;



data[0]=32'b00000000000000000000000000000000;
data[1]=32'b00000000000000000000000000000000;
data[2]=32'b01110000000000000000000000000000;
data[3]=32'b01010001000000000000000000000001;
data[4]=32'b01000001010000100000110000000000;
data[5]=32'b11110010010000000000000000000010;
data[6]=32'b11110010100000000000000000001000;
data[7]=32'b11100001100000100000000000000000;
data[8]=32'b01110001110001100001000000000000;
data[9]=32'b10110000000010100000000000000000;
data[10]=32'b01000001000001100000000000000000;
data[11]=32'b01010000100000100000000000000001;
data[12]=32'b01110001110000100001010000000000;
data[13]=32'b10010000000010010000000000000000;
data[14]=32'b01010001000001000000000000000000;



//data[23] = 32'b00000000000000000000000000000000;
//data[24] = 32'b00000000000000000000000000000000;
//data[25] = 32'b00000000000000000000000000000000;
//data[26] = 32'b00000000000000000000000000000000;
//data[27] = 32'b00000000000000000000000000000000;
//data[28] = 32'b00000000000000000000000000000000;
//data[29] = 32'b00000000000000000000000000000000;
//data[30] = 32'b00000000000000000000000000000000;
//data[31] = 32'b00000000000000000000000000000000;
//data[32] = 32'b00000000000000000000000000000000;
//data[33] = 32'b00000000000000000000000000000000;
//data[34] = 32'b00000000000000000000000000000000;
//data[35] = 32'b00000000000000000000000000000000;
//data[36] = 32'b00000000000000000000000000000000;
//data[37] = 32'b00000000000000000000000000000000;
//data[38] = 32'b00000000000000000000000000000000;
//data[39] = 32'b00000000000000000000000000000000;
//data[40] = 32'b00000000000000000000000000000000;
//data[41] = 32'b00000000000000000000000000000000;
//data[42] = 32'b00000000000000000000000000000000;
//data[43] = 32'b00000000000000000000000000000000;
//data[44] = 32'b00000000000000000000000000000000;
//data[45] = 32'b00000000000000000000000000000000;
//data[46] = 32'b00000000000000000000000000000000;
//data[47] = 32'b00000000000000000000000000000000;
//data[48] = 32'b00000000000000000000000000000000;
//data[49] = 32'b00000000000000000000000000000000;
//data[50] = 32'b00000000000000000000000000000000;
//data[51] = 32'b00000000000000000000000000000000;
//data[52] = 32'b00000000000000000000000000000000;
//data[53] = 32'b00000000000000000000000000000000;
//data[54] = 32'b00000000000000000000000000000000;
//data[55] = 32'b00000000000000000000000000000000;
//data[56] = 32'b00000000000000000000000000000000;
//data[57] = 32'b00000000000000000000000000000000;
//data[58] = 32'b00000000000000000000000000000000;
//data[59] = 32'b00000000000000000000000000000000;
end

always @(posedge clock) begin
insto=data[addr+2];
ip=data[add+1];
idp=data[addr]
end
endmodule