`timescale 1ns / 1ps
`include "ifetch.v"
`include "IF_ID_buffer.v"

module stage1 (
    ports
);
    
endmodule